library Common;
  use Common.CommonLib.all;

ARCHITECTURE studentVersion OF envelopeRetreiver IS
BEGIN

  morseEnvelope <= '0';

END ARCHITECTURE studentVersion;
