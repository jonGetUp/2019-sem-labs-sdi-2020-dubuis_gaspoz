ARCHITECTURE studentVersion OF resizer IS
BEGIN
  resizeOut <= (others => '0');
END ARCHITECTURE studentVersion;
