ARCHITECTURE studentVersion OF parallelAdder IS
BEGIN

  sum <= (others => '0');
  cOut <= '0';

END ARCHITECTURE studentVersion;
