ARCHITECTURE studentVersion OF periphSpeedController IS
BEGIN
  enableOut <= '0';
END ARCHITECTURE studentVersion;
