ARCHITECTURE studentVersion OF characterRegister IS
BEGIN

  charOut <= (others => '0');

END ARCHITECTURE studentVersion;
