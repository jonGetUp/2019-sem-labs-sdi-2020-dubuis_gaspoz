ARCHITECTURE studentVersion OF sawtoothToTriangle IS
BEGIN
  triangle <= (others => '0');
END ARCHITECTURE studentVersion;
