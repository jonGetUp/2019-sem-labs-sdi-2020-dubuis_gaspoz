ARCHITECTURE studentVersion OF periphSizeReg IS
BEGIN
  patternSize <= (others => '0');
END ARCHITECTURE studentVersion;
