ARCHITECTURE studentVersion OF pipelineAdder IS
BEGIN

  sum <= (others => '0');
  cOut <= '0';

END ARCHITECTURE studentVersion;
