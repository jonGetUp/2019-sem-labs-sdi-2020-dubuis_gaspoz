ARCHITECTURE studentVersion OF interpolatorCalculatePolynom IS
BEGIN
  sampleOut <= (others => '0');
END ARCHITECTURE studentVersion;
