ARCHITECTURE order2_studentVersion OF DAC IS
BEGIN
  serialOut <= '0';
END ARCHITECTURE order2_studentVersion;
