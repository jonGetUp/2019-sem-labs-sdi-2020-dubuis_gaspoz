ARCHITECTURE studentVersion OF interpolatorCoefficients IS
BEGIN
  a <= (others => '0');
  b <= (others => '0');
  c <= (others => '0');
  d <= (others => '0');
END ARCHITECTURE studentVersion;
