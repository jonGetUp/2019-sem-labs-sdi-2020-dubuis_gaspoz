LIBRARY ieee;
  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;

PACKAGE beamerTest_pck IS

  function trim_X (arg : signed) return signed;

END beamerTest_pck;
