ARCHITECTURE studentVersion OF morseToCharDecoder IS
BEGIN

  charValid <= '0';
  charOut <= (others => '0');

END ARCHITECTURE studentVersion;
