ARCHITECTURE studentVersion OF interpolatorShiftRegister IS
BEGIN
  sample1 <= (others => '0');
  sample2 <= (others => '0');
  sample3 <= (others => '0');
  sample4 <= (others => '0');
END ARCHITECTURE studentVersion;
