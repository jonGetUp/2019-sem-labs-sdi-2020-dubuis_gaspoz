ARCHITECTURE studentVersion OF periphAddressDecoder IS
BEGIN
  selControl  <= '0';
--  selSize     <= '0';
  selSpeed    <= '0';
  selX        <= '0';
  selY        <= '0';
  selZ        <= '0';
END ARCHITECTURE studentVersion;

