ARCHITECTURE studentVersion OF sinCosTable IS
BEGIN
  sine <= (others => '0');
  cosine <= (others => '0');
END ARCHITECTURE studentVersion;
