ARCHITECTURE studentVersion OF blockRAMAddressCounter IS
BEGIN
  addr <= (others => '0');
END ARCHITECTURE studentVersion;
