ARCHITECTURE studentVersion OF sawtoothGen IS
BEGIN
  sawtooth <= (others => '0');
END ARCHITECTURE studentVersion;

