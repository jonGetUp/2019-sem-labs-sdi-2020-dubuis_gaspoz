ARCHITECTURE studentVersion OF offsetToUnsigned IS
BEGIN
  unsignedOut <= (others => '0');
END ARCHITECTURE studentVersion;
