ARCHITECTURE studentVersion OF blockRAMControl IS
BEGIN
  cntIncr <= '0';
  memWr   <= '0';
  memEn   <= '0';
END ARCHITECTURE studentVersion;
