ARCHITECTURE studentVersion OF triangleToPolygon IS
BEGIN
  polygon <= (others => '0');
END ARCHITECTURE studentVersion;
