ARCHITECTURE studentVersion OF sawtoothToSquare IS
BEGIN
  square <= (others => '0');
END ARCHITECTURE studentVersion;
