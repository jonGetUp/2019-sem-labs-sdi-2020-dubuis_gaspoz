ARCHITECTURE studentVersion OF DAC IS
BEGIN
  serialOut <= '0';
END ARCHITECTURE studentVersion;
