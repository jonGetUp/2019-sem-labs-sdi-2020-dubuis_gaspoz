ARCHITECTURE studentVersion OF interpolatorTrigger IS
BEGIN
  triggerOut <= '0';
END ARCHITECTURE studentVersion;
