ARCHITECTURE studentVersion OF periphControlReg IS
BEGIN
  run               <= '0';
  updatePattern     <= '0';
  interpolateLinear <= '0';
END ARCHITECTURE studentVersion;
