ARCHITECTURE studentVersion OF periphSpeedReg IS
BEGIN
  updatePeriod <= (others => '0');
END ARCHITECTURE studentVersion;

