ARCHITECTURE studentVersion OF lowpass IS
BEGIN
  lowpassOut <= (others => '0');
END ARCHITECTURE studentVersion;
